* Current Mirror Netlist
M1 out in VDD VDD PMOS L=0.18u W=10u
M2 in in VDD VDD PMOS L=0.18u W=10u
R1 out VDD 1k
.END
